module fetch_seq(
   
